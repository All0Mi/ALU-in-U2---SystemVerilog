`ifndef ALU_DEF

`define ALU_DEF
`include "./bit_set/bit_set.sv"
`include "./bit_shift/bit_shift.sv"
`include "./comparator/comparator.sv"
`include "./u2_to_sm/u2_to_sm.sv"
`include "./MUX.sv"
`include "./reg.sv"
  
`endif